module OR_Gate(
    input1,
    input2,
    result
);

input	input1, input2;
output	result;

assign result = input1 | input2;

endmodule
